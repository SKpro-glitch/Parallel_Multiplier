// -----------------------------------------------------------------------------
// Copyright 2024 Soham Kapur
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
// Project Name: Parameterized Parallel Multiplier
// Description:  This module creates a combinational intermediate product for the Wallace Tree multiplier, which is one stage of the Carry Save Adder.
// -----------------------------------------------------------------------------

`timescale 1ns / 1ps

//Intermediate product calculation
module Inter_Prod #(parameter bits = 31)(
    input [bits:0] x, y, z,
    output [bits:0] s, c
    );
    
    //Combinational Implementation of Full Adder
    assign s = x ^ y ^ z;
    assign c = (x & y) | (y & z) | (x & z);
    
endmodule
